
`ifndef TEMPLATE_MASTER_SEQUENCER_SV
`define TEMPLATE_MASTER_SEQUENCER_SV

function template_master_sequencer::new (string name, uvm_component parent);
  super.new(name, parent);
endfunction : new

`endif // TEMPLATE_MASTER_SEQUENCER_SV


