
`ifndef TEMPLATE_PKG_SV
`define TEMPLATE_PKG_SV

package template_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "template.svh"

endpackage : template_pkg

   
`endif //  `ifndef TEMPLATE_PKG_SV
